LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FULL_COLOR_LED IS
PORT(
	RESETN, CLK : IN STD_LOGIC;
	
	R_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	G_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	B_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	R : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	G : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	B : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END FULL_COLOR_LED;

ARCHITECTURE HB OF FULL_COLOR_LED IS

SIGNAL CNT : INTEGER RANGE 0 TO 100;

SIGNAL R_REG : INTEGER RANGE 0 TO 100;
SIGNAL G_REG : INTEGER RANGE 0 TO 100;
SIGNAL B_REG : INTEGER RANGE 0 TO 100;

BEGIN

-- SWITCH REG

PROCESS(RESETN, CLK)
BEGIN	
	IF RESETN = '1' THEN
		R_REG <= 0;
		G_REG <= 0;
		B_REG <= 0;
	ELSIF CLK'EVENT AND CLK = '1' THEN
		CASE R_IN IS
			WHEN "0001" => R_REG <= 0;   -- DUTY 0%
			WHEN "0010" => R_REG <= 33;-- DUTY 33%
			WHEN "0100" => R_REG <= 66;-- DUTY 66%
			WHEN "1000" => R_REG <= 100;-- DUTY 100%
			WHEN OTHERS => NULL;
		END CASE;
		
		CASE G_IN IS
			WHEN "0001" => G_REG <= 0;   -- DUTY 0%
			WHEN "0010" => G_REG <= 33;-- DUTY 33%
			WHEN "0100" => G_REG <= 66;-- DUTY 66%
			WHEN "1000" => G_REG <= 100;-- DUTY 100%
			WHEN OTHERS => NULL;
		END CASE;

		CASE B_IN IS
			WHEN "0001" => B_REG <= 0;   -- DUTY 0%
			WHEN "0010" => B_REG <= 33;-- DUTY 33%
			WHEN "0100" => B_REG <= 66;-- DUTY 66%
			WHEN "1000" => B_REG <= 100;-- DUTY 100%
			WHEN OTHERS => NULL;
		END CASE;
	END IF;
END PROCESS;
		
PROCESS(RESETN, CLK)
BEGIN	
	IF RESETN = '1' THEN
		CNT <= 0;
	ELSIF CLK'EVENT AND CLK = '1' THEN
		IF CNT >= 99 THEN	
			CNT <= 0;
		ELSE
			CNT <= CNT + 1;
		END IF;
	END IF;
END PROCESS;

R <= "1111" WHEN CNT < R_REG ELSE "0000";
G <= "1111" WHEN CNT < G_REG ELSE "0000";
B <= "1111" WHEN CNT < B_REG ELSE "0000";

END HB;

			

	
